`line 4
module vloga_dig_submod_conso_dyn_bd(capa_charge_val,internal_energy,fin_test,\_ana_evt_sig_#1#66#\ ,\_ana_evt_sig_#2#69#\ );
parameter real alim_voltage = 0.0;
parameter real slew_lower_threshold_pct = 0.0;
parameter real slew_upper_threshold_pct = 0.0;
parameter real input_threshold_pct = 0.0;
parameter real output_threshold_pct = 0.0;
input wreal capa_charge_val ;
output wreal internal_energy ;
input  fin_test ;
input  \_ana_evt_sig_#1#66#\  ;
input  \_ana_evt_sig_#2#69#\  ;
endmodule

