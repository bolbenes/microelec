`line 4
module vloga_dig_submod_input_capa_bd(capa_charge_val,capa_test_val,circuit_propagation_time,test_propagation_time,fin_test,\_ana_evt_sig_#1#73#\ ,\_ana_evt_sig_#2#76#\ ,\_ana_evt_sig_#3#79#\ ,\_ana_evt_sig_#4#82#\ ,\_ana_evt_sig_#5#85#\ ,\_ana_evt_sig_#6#88#\ );
parameter real alim_voltage = 0.0;
parameter real slew_lower_threshold_pct = 0.0;
parameter real slew_upper_threshold_pct = 0.0;
parameter real input_threshold_pct = 0.0;
parameter real output_threshold_pct = 0.0;
input wreal capa_charge_val ;
input wreal capa_test_val ;
output wreal circuit_propagation_time ;
output wreal test_propagation_time ;
input  fin_test ;
input  \_ana_evt_sig_#1#73#\  ;
input  \_ana_evt_sig_#2#76#\  ;
input  \_ana_evt_sig_#3#79#\  ;
input  \_ana_evt_sig_#4#82#\  ;
input  \_ana_evt_sig_#5#85#\  ;
input  \_ana_evt_sig_#6#88#\  ;
endmodule

