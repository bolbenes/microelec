LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

LIBRARY STD;
USE STD.ALL;

ENTITY cmos_transition IS
  GENERIC (
   alpha_threshold :   real :=  2.176097e+01;
   slew_lower_threshold_pct :   real :=  3.000000e-01;
   slew_upper_threshold_pct :   real :=  7.000000e-01;
   tt_tablex :   real_vector(0 to 478) := ( 0.000000e+00 , 1.987305e-01 , 2.270508e-01 , 2.443848e-01 , 2.573242e-01 , 2.678223e-01 , 2.766113e-01 , 2.844238e-01 , 2.912598e-01 , 2.976074e-01 , 3.032227e-01 , 3.085938e-01 , 3.134766e-01 , 3.181152e-01 , 3.225098e-01 , 3.266602e-01 , 3.305664e-01 , 3.344727e-01 , 3.381348e-01 , 3.417969e-01 , 3.452148e-01 , 3.483887e-01 , 3.515625e-01 , 3.547363e-01 , 3.576660e-01 , 3.605957e-01 , 3.635254e-01 , 3.662109e-01 , 3.688965e-01 , 3.715820e-01 , 3.740234e-01 , 3.764648e-01 , 3.789062e-01 , 3.813477e-01 , 3.835449e-01 , 3.857422e-01 , 3.879395e-01 , 3.901367e-01 , 3.923340e-01 , 3.945312e-01 , 3.964844e-01 , 3.984375e-01 , 4.003906e-01 , 4.023438e-01 , 4.042969e-01 , 4.062500e-01 , 4.079590e-01 , 4.096680e-01 , 4.113770e-01 , 4.130859e-01 , 4.147949e-01 , 4.165039e-01 , 4.182129e-01 , 4.199219e-01 , 4.213867e-01 , 4.228516e-01 , 4.243164e-01 , 4.257812e-01 , 4.272461e-01 , 4.287109e-01 , 4.301758e-01 , 4.316406e-01 , 4.331055e-01 , 4.345703e-01 , 4.357910e-01 , 4.370117e-01 , 4.382324e-01 , 4.394531e-01 , 4.406738e-01 , 4.418945e-01 , 4.431152e-01 , 4.443359e-01 , 4.455566e-01 , 4.467773e-01 , 4.479980e-01 , 4.492188e-01 , 4.501953e-01 , 4.511719e-01 , 4.521484e-01 , 4.531250e-01 , 4.541016e-01 , 4.550781e-01 , 4.560547e-01 , 4.570312e-01 , 4.580078e-01 , 4.589844e-01 , 4.599609e-01 , 4.609375e-01 , 4.619141e-01 , 4.628906e-01 , 4.638672e-01 , 4.648438e-01 , 4.655762e-01 , 4.663086e-01 , 4.670410e-01 , 4.677734e-01 , 4.685059e-01 , 4.692383e-01 , 4.699707e-01 , 4.707031e-01 , 4.714355e-01 , 4.721680e-01 , 4.729004e-01 , 4.736328e-01 , 4.743652e-01 , 4.750977e-01 , 4.758301e-01 , 4.765625e-01 , 4.772949e-01 , 4.780273e-01 , 4.787598e-01 , 4.792480e-01 , 4.797363e-01 , 4.802246e-01 , 4.807129e-01 , 4.812012e-01 , 4.816895e-01 , 4.821777e-01 , 4.826660e-01 , 4.831543e-01 , 4.836426e-01 , 4.841309e-01 , 4.846191e-01 , 4.851074e-01 , 4.855957e-01 , 4.860840e-01 , 4.865723e-01 , 4.870605e-01 , 4.875488e-01 , 4.880371e-01 , 4.885254e-01 , 4.890137e-01 , 4.895020e-01 , 4.899902e-01 , 4.904785e-01 , 4.909668e-01 , 4.914551e-01 , 4.919434e-01 , 4.921875e-01 , 4.924316e-01 , 4.926758e-01 , 4.929199e-01 , 4.931641e-01 , 4.934082e-01 , 4.936523e-01 , 4.938965e-01 , 4.941406e-01 , 4.943848e-01 , 4.946289e-01 , 4.948730e-01 , 4.951172e-01 , 4.953613e-01 , 4.956055e-01 , 4.958496e-01 , 4.960938e-01 , 4.963379e-01 , 4.965820e-01 , 4.968262e-01 , 4.970703e-01 , 4.973145e-01 , 4.975586e-01 , 4.978027e-01 , 4.980469e-01 , 4.982910e-01 , 4.985352e-01 , 4.987793e-01 , 4.990234e-01 , 4.992676e-01 , 4.995117e-01 , 4.997559e-01 , 5.000000e-01 , 5.002441e-01 , 5.004883e-01 , 5.007324e-01 , 5.009766e-01 , 5.012207e-01 , 5.014648e-01 , 5.017090e-01 , 5.019531e-01 , 5.021973e-01 , 5.024414e-01 , 5.026856e-01 , 5.029297e-01 , 5.031738e-01 , 5.034180e-01 , 5.036621e-01 , 5.039062e-01 , 5.041504e-01 , 5.043945e-01 , 5.046387e-01 , 5.048828e-01 , 5.051269e-01 , 5.053711e-01 , 5.056152e-01 , 5.058594e-01 , 5.061035e-01 , 5.063477e-01 , 5.065918e-01 , 5.068359e-01 , 5.070801e-01 , 5.073242e-01 , 5.075684e-01 , 5.078125e-01 , 5.080566e-01 , 5.083008e-01 , 5.085449e-01 , 5.087891e-01 , 5.090332e-01 , 5.092773e-01 , 5.095215e-01 , 5.097656e-01 , 5.100098e-01 , 5.102539e-01 , 5.104981e-01 , 5.107422e-01 , 5.109863e-01 , 5.112305e-01 , 5.114746e-01 , 5.117188e-01 , 5.119629e-01 , 5.122070e-01 , 5.124512e-01 , 5.126953e-01 , 5.129394e-01 , 5.131836e-01 , 5.134277e-01 , 5.136719e-01 , 5.139160e-01 , 5.141602e-01 , 5.144043e-01 , 5.146484e-01 , 5.148926e-01 , 5.151367e-01 , 5.153809e-01 , 5.156250e-01 , 5.158691e-01 , 5.161133e-01 , 5.163574e-01 , 5.166016e-01 , 5.168457e-01 , 5.170898e-01 , 5.173340e-01 , 5.175781e-01 , 5.178223e-01 , 5.180664e-01 , 5.183106e-01 , 5.185547e-01 , 5.187988e-01 , 5.190430e-01 , 5.192871e-01 , 5.195312e-01 , 5.197754e-01 , 5.200195e-01 , 5.202637e-01 , 5.205078e-01 , 5.207519e-01 , 5.209961e-01 , 5.212402e-01 , 5.214844e-01 , 5.217285e-01 , 5.219727e-01 , 5.222168e-01 , 5.224609e-01 , 5.227051e-01 , 5.229492e-01 , 5.231934e-01 , 5.234375e-01 , 5.236816e-01 , 5.239258e-01 , 5.241699e-01 , 5.244141e-01 , 5.246582e-01 , 5.249023e-01 , 5.251465e-01 , 5.253906e-01 , 5.256348e-01 , 5.258789e-01 , 5.261231e-01 , 5.263672e-01 , 5.266113e-01 , 5.268555e-01 , 5.270996e-01 , 5.273438e-01 , 5.275879e-01 , 5.278320e-01 , 5.280762e-01 , 5.283203e-01 , 5.285644e-01 , 5.288086e-01 , 5.290527e-01 , 5.292969e-01 , 5.295410e-01 , 5.297852e-01 , 5.300293e-01 , 5.302734e-01 , 5.305176e-01 , 5.307617e-01 , 5.310059e-01 , 5.312500e-01 , 5.314941e-01 , 5.317383e-01 , 5.319824e-01 , 5.322266e-01 , 5.324707e-01 , 5.327148e-01 , 5.329590e-01 , 5.332031e-01 , 5.334473e-01 , 5.336914e-01 , 5.339356e-01 , 5.341797e-01 , 5.344238e-01 , 5.346680e-01 , 5.349121e-01 , 5.351562e-01 , 5.354004e-01 , 5.356445e-01 , 5.358887e-01 , 5.361328e-01 , 5.363769e-01 , 5.366211e-01 , 5.368652e-01 , 5.371094e-01 , 5.373535e-01 , 5.375977e-01 , 5.378418e-01 , 5.380859e-01 , 5.383301e-01 , 5.385742e-01 , 5.388184e-01 , 5.390625e-01 , 5.393066e-01 , 5.395508e-01 , 5.400391e-01 , 5.405273e-01 , 5.410156e-01 , 5.415039e-01 , 5.419922e-01 , 5.424805e-01 , 5.429688e-01 , 5.434570e-01 , 5.439453e-01 , 5.444336e-01 , 5.449219e-01 , 5.454102e-01 , 5.458984e-01 , 5.463867e-01 , 5.468750e-01 , 5.473633e-01 , 5.478516e-01 , 5.483398e-01 , 5.488281e-01 , 5.493164e-01 , 5.498047e-01 , 5.502930e-01 , 5.507812e-01 , 5.512695e-01 , 5.517578e-01 , 5.522461e-01 , 5.527344e-01 , 5.532227e-01 , 5.537109e-01 , 5.541992e-01 , 5.546875e-01 , 5.551758e-01 , 5.556641e-01 , 5.561523e-01 , 5.566406e-01 , 5.571289e-01 , 5.578613e-01 , 5.585938e-01 , 5.593262e-01 , 5.600586e-01 , 5.607910e-01 , 5.615234e-01 , 5.622559e-01 , 5.629883e-01 , 5.637207e-01 , 5.644531e-01 , 5.651856e-01 , 5.659180e-01 , 5.666504e-01 , 5.673828e-01 , 5.681152e-01 , 5.688477e-01 , 5.695801e-01 , 5.703125e-01 , 5.710449e-01 , 5.717773e-01 , 5.725098e-01 , 5.732422e-01 , 5.739746e-01 , 5.747070e-01 , 5.754394e-01 , 5.761719e-01 , 5.771484e-01 , 5.781250e-01 , 5.791016e-01 , 5.800781e-01 , 5.810547e-01 , 5.820312e-01 , 5.830078e-01 , 5.839844e-01 , 5.849609e-01 , 5.859375e-01 , 5.869141e-01 , 5.878906e-01 , 5.888672e-01 , 5.898438e-01 , 5.908203e-01 , 5.917969e-01 , 5.927734e-01 , 5.937500e-01 , 5.949707e-01 , 5.961914e-01 , 5.974121e-01 , 5.986328e-01 , 5.998535e-01 , 6.010742e-01 , 6.022949e-01 , 6.035156e-01 , 6.047363e-01 , 6.059570e-01 , 6.071777e-01 , 6.083984e-01 , 6.096191e-01 , 6.110840e-01 , 6.125488e-01 , 6.140137e-01 , 6.154785e-01 , 6.169434e-01 , 6.184082e-01 , 6.198731e-01 , 6.213379e-01 , 6.228027e-01 , 6.242676e-01 , 6.259766e-01 , 6.276856e-01 , 6.293945e-01 , 6.311035e-01 , 6.328125e-01 , 6.345215e-01 , 6.362305e-01 , 6.381836e-01 , 6.401367e-01 , 6.420898e-01 , 6.440430e-01 , 6.459961e-01 , 6.479492e-01 , 6.501465e-01 , 6.523438e-01 , 6.545410e-01 , 6.567383e-01 , 6.591797e-01 , 6.616211e-01 , 6.640625e-01 , 6.667481e-01 , 6.694336e-01 , 6.721191e-01 , 6.750488e-01 , 6.779785e-01 , 6.811523e-01 , 6.845703e-01 , 6.879883e-01 , 6.916504e-01 , 6.955566e-01 , 6.997070e-01 , 7.041016e-01 , 7.089844e-01 , 7.141113e-01 , 7.197266e-01 , 7.260742e-01 , 7.331543e-01 , 7.414551e-01 , 7.514648e-01 , 7.641602e-01 , 7.817383e-01 , 8.122559e-01 , 1.000000e+00 ) ;
   tt_tabley :   real_vector(0 to 478) := ( 0.000000e+00 , 1.004040e-03 , 2.011870e-03 , 3.015290e-03 , 4.025590e-03 , 5.046610e-03 , 6.057610e-03 , 7.087980e-03 , 8.100070e-03 , 9.138600e-03 , 1.014055e-02 , 1.117319e-02 , 1.218047e-02 , 1.319657e-02 , 1.421583e-02 , 1.523114e-02 , 1.623378e-02 , 1.728333e-02 , 1.831201e-02 , 1.938175e-02 , 2.042108e-02 , 2.142259e-02 , 2.245653e-02 , 2.352825e-02 , 2.454866e-02 , 2.560066e-02 , 2.668498e-02 , 2.770682e-02 , 2.875938e-02 , 2.983871e-02 , 3.084680e-02 , 3.188008e-02 , 3.293915e-02 , 3.402535e-02 , 3.502547e-02 , 3.604809e-02 , 3.709377e-02 , 3.816234e-02 , 3.925593e-02 , 4.037449e-02 , 4.139030e-02 , 4.242694e-02 , 4.348497e-02 , 4.456499e-02 , 4.566765e-02 , 4.679362e-02 , 4.779853e-02 , 4.882235e-02 , 4.986562e-02 , 5.092891e-02 , 5.201283e-02 , 5.311801e-02 , 5.424513e-02 , 5.539492e-02 , 5.639906e-02 , 5.742092e-02 , 5.846103e-02 , 5.951996e-02 , 6.059831e-02 , 6.169670e-02 , 6.281582e-02 , 6.395636e-02 , 6.511907e-02 , 6.630474e-02 , 6.731094e-02 , 6.833421e-02 , 6.937509e-02 , 7.043418e-02 , 7.151203e-02 , 7.260931e-02 , 7.372667e-02 , 7.486496e-02 , 7.602472e-02 , 7.720696e-02 , 7.841247e-02 , 7.964217e-02 , 8.064401e-02 , 8.166249e-02 , 8.269822e-02 , 8.375170e-02 , 8.482360e-02 , 8.591459e-02 , 8.702537e-02 , 8.815667e-02 , 8.930930e-02 , 9.048410e-02 , 9.168195e-02 , 9.290382e-02 , 9.415076e-02 , 9.542377e-02 , 9.672414e-02 , 9.805305e-02 , 9.906939e-02 , 1.001031e-01 , 1.011546e-01 , 1.022253e-01 , 1.033152e-01 , 1.044255e-01 , 1.055567e-01 , 1.067100e-01 , 1.078861e-01 , 1.090862e-01 , 1.103114e-01 , 1.115624e-01 , 1.128409e-01 , 1.141482e-01 , 1.154854e-01 , 1.168544e-01 , 1.182567e-01 , 1.196940e-01 , 1.211686e-01 , 1.221734e-01 , 1.231963e-01 , 1.242381e-01 , 1.252996e-01 , 1.263817e-01 , 1.274850e-01 , 1.286108e-01 , 1.297600e-01 , 1.309336e-01 , 1.321327e-01 , 1.333588e-01 , 1.346131e-01 , 1.358971e-01 , 1.372115e-01 , 1.385605e-01 , 1.399434e-01 , 1.413632e-01 , 1.428220e-01 , 1.443221e-01 , 1.458662e-01 , 1.474571e-01 , 1.490980e-01 , 1.507921e-01 , 1.525434e-01 , 1.543560e-01 , 1.562347e-01 , 1.581841e-01 , 1.591872e-01 , 1.602102e-01 , 1.612540e-01 , 1.623193e-01 , 1.634070e-01 , 1.645183e-01 , 1.656539e-01 , 1.668150e-01 , 1.680028e-01 , 1.692183e-01 , 1.704630e-01 , 1.717380e-01 , 1.730447e-01 , 1.743848e-01 , 1.757597e-01 , 1.771710e-01 , 1.786206e-01 , 1.801103e-01 , 1.816420e-01 , 1.832178e-01 , 1.848399e-01 , 1.865104e-01 , 1.882317e-01 , 1.900064e-01 , 1.918371e-01 , 1.937264e-01 , 1.956771e-01 , 1.976921e-01 , 1.997744e-01 , 2.019271e-01 , 2.041532e-01 , 2.064559e-01 , 2.088383e-01 , 2.113036e-01 , 2.138550e-01 , 2.164953e-01 , 2.192276e-01 , 2.220546e-01 , 2.249788e-01 , 2.280026e-01 , 2.311280e-01 , 2.343568e-01 , 2.376903e-01 , 2.411296e-01 , 2.446751e-01 , 2.483271e-01 , 2.520852e-01 , 2.559487e-01 , 2.599165e-01 , 2.639869e-01 , 2.681581e-01 , 2.724276e-01 , 2.767927e-01 , 2.812506e-01 , 2.857981e-01 , 2.904317e-01 , 2.951479e-01 , 2.999432e-01 , 3.048136e-01 , 3.097556e-01 , 3.147653e-01 , 3.198391e-01 , 3.249725e-01 , 3.301634e-01 , 3.354073e-01 , 3.407011e-01 , 3.460412e-01 , 3.514247e-01 , 3.568483e-01 , 3.623091e-01 , 3.678043e-01 , 3.733312e-01 , 3.788872e-01 , 3.844698e-01 , 3.900766e-01 , 3.957054e-01 , 4.013539e-01 , 4.070202e-01 , 4.127022e-01 , 4.183981e-01 , 4.241059e-01 , 4.298239e-01 , 4.355505e-01 , 4.412839e-01 , 4.470226e-01 , 4.527649e-01 , 4.585095e-01 , 4.642548e-01 , 4.699994e-01 , 4.757418e-01 , 4.814807e-01 , 4.872146e-01 , 4.929421e-01 , 4.986620e-01 , 5.043728e-01 , 5.100731e-01 , 5.157616e-01 , 5.214369e-01 , 5.270976e-01 , 5.327423e-01 , 5.383695e-01 , 5.439778e-01 , 5.495657e-01 , 5.551317e-01 , 5.606743e-01 , 5.661918e-01 , 5.716826e-01 , 5.771451e-01 , 5.825777e-01 , 5.879784e-01 , 5.933456e-01 , 5.986774e-01 , 6.039719e-01 , 6.092271e-01 , 6.144412e-01 , 6.196119e-01 , 6.247374e-01 , 6.298153e-01 , 6.348437e-01 , 6.398202e-01 , 6.447426e-01 , 6.496087e-01 , 6.544162e-01 , 6.591629e-01 , 6.638464e-01 , 6.684646e-01 , 6.730152e-01 , 6.774961e-01 , 6.819051e-01 , 6.862402e-01 , 6.904995e-01 , 6.946813e-01 , 6.987838e-01 , 7.028055e-01 , 7.067452e-01 , 7.106016e-01 , 7.143738e-01 , 7.180611e-01 , 7.216630e-01 , 7.251792e-01 , 7.286097e-01 , 7.319547e-01 , 7.352146e-01 , 7.383901e-01 , 7.414820e-01 , 7.444915e-01 , 7.474197e-01 , 7.502682e-01 , 7.530386e-01 , 7.557325e-01 , 7.583519e-01 , 7.608987e-01 , 7.633749e-01 , 7.657826e-01 , 7.681239e-01 , 7.704010e-01 , 7.726161e-01 , 7.747713e-01 , 7.768687e-01 , 7.789105e-01 , 7.808987e-01 , 7.828354e-01 , 7.847225e-01 , 7.865621e-01 , 7.883558e-01 , 7.901056e-01 , 7.918133e-01 , 7.934804e-01 , 7.951086e-01 , 7.966994e-01 , 7.982543e-01 , 7.997748e-01 , 8.012622e-01 , 8.027178e-01 , 8.041429e-01 , 8.055385e-01 , 8.069060e-01 , 8.082462e-01 , 8.095605e-01 , 8.108494e-01 , 8.121140e-01 , 8.133554e-01 , 8.145742e-01 , 8.157714e-01 , 8.169476e-01 , 8.181037e-01 , 8.192402e-01 , 8.203580e-01 , 8.214575e-01 , 8.225394e-01 , 8.236044e-01 , 8.246528e-01 , 8.256854e-01 , 8.267025e-01 , 8.277047e-01 , 8.296660e-01 , 8.315727e-01 , 8.334282e-01 , 8.352351e-01 , 8.369962e-01 , 8.387140e-01 , 8.403907e-01 , 8.420283e-01 , 8.436289e-01 , 8.451941e-01 , 8.467258e-01 , 8.482253e-01 , 8.496942e-01 , 8.511337e-01 , 8.525452e-01 , 8.539298e-01 , 8.552885e-01 , 8.566225e-01 , 8.579327e-01 , 8.592200e-01 , 8.604852e-01 , 8.617292e-01 , 8.629527e-01 , 8.641564e-01 , 8.653410e-01 , 8.665072e-01 , 8.676555e-01 , 8.687866e-01 , 8.699009e-01 , 8.709990e-01 , 8.720814e-01 , 8.731485e-01 , 8.742009e-01 , 8.752389e-01 , 8.762629e-01 , 8.772734e-01 , 8.787644e-01 , 8.802270e-01 , 8.816621e-01 , 8.830709e-01 , 8.844543e-01 , 8.858132e-01 , 8.871486e-01 , 8.884612e-01 , 8.897518e-01 , 8.910211e-01 , 8.922699e-01 , 8.934987e-01 , 8.947083e-01 , 8.958991e-01 , 8.970718e-01 , 8.982269e-01 , 8.993650e-01 , 9.004864e-01 , 9.015917e-01 , 9.026812e-01 , 9.037555e-01 , 9.048149e-01 , 9.058598e-01 , 9.068905e-01 , 9.079075e-01 , 9.089111e-01 , 9.102289e-01 , 9.115240e-01 , 9.127974e-01 , 9.140495e-01 , 9.152810e-01 , 9.164925e-01 , 9.176847e-01 , 9.188579e-01 , 9.200128e-01 , 9.211499e-01 , 9.222695e-01 , 9.233722e-01 , 9.244584e-01 , 9.255284e-01 , 9.265828e-01 , 9.276218e-01 , 9.286458e-01 , 9.296552e-01 , 9.308968e-01 , 9.321167e-01 , 9.333155e-01 , 9.344937e-01 , 9.356519e-01 , 9.367905e-01 , 9.379100e-01 , 9.390110e-01 , 9.400938e-01 , 9.411589e-01 , 9.422067e-01 , 9.432375e-01 , 9.442518e-01 , 9.454476e-01 , 9.466207e-01 , 9.477716e-01 , 9.489008e-01 , 9.500089e-01 , 9.510963e-01 , 9.521635e-01 , 9.532110e-01 , 9.542392e-01 , 9.552485e-01 , 9.564025e-01 , 9.575320e-01 , 9.586374e-01 , 9.597192e-01 , 9.607781e-01 , 9.618144e-01 , 9.628286e-01 , 9.639613e-01 , 9.650664e-01 , 9.661446e-01 , 9.671963e-01 , 9.682223e-01 , 9.692229e-01 , 9.703190e-01 , 9.713845e-01 , 9.724200e-01 , 9.734261e-01 , 9.745105e-01 , 9.755602e-01 , 9.765761e-01 , 9.776554e-01 , 9.786958e-01 , 9.796982e-01 , 9.807494e-01 , 9.817577e-01 , 9.828029e-01 , 9.838752e-01 , 9.848936e-01 , 9.859269e-01 , 9.869653e-01 , 9.879997e-01 , 9.890207e-01 , 9.900701e-01 , 9.910808e-01 , 9.920871e-01 , 9.931070e-01 , 9.941091e-01 , 9.951203e-01 , 9.961331e-01 , 9.971441e-01 , 9.981473e-01 , 9.991521e-01 , 1.000000e+00 )  );
  PORT (
    SIGNAL din : IN STD_LOGIC;
    SIGNAL dout : OUT STD_LOGIC;
    SIGNAL tt_val : IN real);
END ENTITY cmos_transition;

