`line 4
module vloga_dig_submod_input_capa_bd(capa_charge_val,capa_test_val,circuit_propagation_time,test_propagation_time,fin_test,\_ana_evt_sig_#1#74#\ ,\_ana_evt_sig_#2#77#\ ,\_ana_evt_sig_#3#80#\ );
parameter real alim_voltage = 0.0;
parameter real slew_lower_threshold_pct = 0.0;
parameter real slew_upper_threshold_pct = 0.0;
parameter real input_threshold_pct = 0.0;
parameter real output_threshold_pct = 0.0;
input wreal capa_charge_val ;
input wreal capa_test_val ;
output wreal circuit_propagation_time ;
output wreal test_propagation_time ;
input  fin_test ;
input  \_ana_evt_sig_#1#74#\  ;
input  \_ana_evt_sig_#2#77#\  ;
input  \_ana_evt_sig_#3#80#\  ;
endmodule

