`line 4
module vloga_dig_submod_hold_study_bd(capa_charge_val,clk_rise_time,d_fall_time,fin_test,\_ana_evt_sig_#1#79#\ ,\_ana_evt_sig_#2#84#\ );
parameter real alim_voltage = 0.0;
parameter real slew_lower_threshold_pct = 0.0;
parameter real slew_upper_threshold_pct = 0.0;
parameter real input_threshold_pct = 0.0;
parameter real output_threshold_pct = 0.0;
input wreal capa_charge_val ;
output wreal clk_rise_time ;
output wreal d_fall_time ;
input  fin_test ;
input  \_ana_evt_sig_#1#79#\  ;
input  \_ana_evt_sig_#2#84#\  ;
endmodule

